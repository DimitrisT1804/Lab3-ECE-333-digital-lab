module VRAM(cord_x, cord_y, colors);
input cord_x, cord_y;
output [2:0] colors;

BRAM_SINGLE_MACRO_RED_inst()

endmodule